`timescale 1ns / 1ps

module cpu_integration_tests_harness ();

  // verilator lint_off PINMISSING
  cpu cpu ();
  // verilator lint_on  PINMISSING
endmodule
