`include "../cpu_core_params.vh"

`ifndef MEMORY_PARAMS_VH
`define MEMORY_PARAMS_VH

// Load/Store types
parameter [LS_SEL_WIDTH:0] LS_TYPE_LOAD_WORD = 0;
parameter [LS_SEL_WIDTH:0] LS_TYPE_LOAD_HALF = 1;
parameter [LS_SEL_WIDTH:0] LS_TYPE_LOAD_HALF_UNSIGNED = 2;
parameter [LS_SEL_WIDTH:0] LS_TYPE_LOAD_BYTE = 3;
parameter [LS_SEL_WIDTH:0] LS_TYPE_LOAD_BYTE_UNSIGNED = 4;
parameter [LS_SEL_WIDTH:0] LS_TYPE_STORE_WORD = 5;
parameter [LS_SEL_WIDTH:0] LS_TYPE_STORE_HALF = 6;
parameter [LS_SEL_WIDTH:0] LS_TYPE_STORE_BYTE = 7;
parameter [LS_SEL_WIDTH:0] LS_TYPE_NONE = 8;

parameter [MEMORY_STATE_WIDTH:0] IDLE = 3'b000;
parameter [MEMORY_STATE_WIDTH:0] READ_SUBMITTING = 3'b001;
parameter [MEMORY_STATE_WIDTH:0] READ_AWAITING = 3'b010;
parameter [MEMORY_STATE_WIDTH:0] READ_SUCCESS = 3'b011;
parameter [MEMORY_STATE_WIDTH:0] WRITE_SUBMITTING = 3'b100;
parameter [MEMORY_STATE_WIDTH:0] WRITE_AWAITING = 3'b101;
parameter [MEMORY_STATE_WIDTH:0] WRITE_SUCCESS = 3'b110;


`endif  // MEMORY_PARAMS_VH
